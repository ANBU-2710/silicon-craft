module uart_top;
endmodule
