module uart_rx;
endmodu
