module clk_div_tb;
endmodule
